// main testbench related parameters 
`define INSTRUCTIONS_FILE "../../main/tb/instructions.txt"
`define RANDOM_DATA_FILE "../../main/tb/random_data.txt"
`define NUMBER_OF_INSTRUCTIONS 10

// clock period
`define T_clk 20
`define half_T_clk 10
// main testbench related parameters 
`define INSTRUCTIONS_FILE "../../main/tb/hex_mc/1-instr_list_no_jump.riscv"
`define DATA_FILE "../../main/tb/hex_mc/min_calc_mem_init.txt"
`define NUMBER_OF_INSTRUCTIONS 10

// clock period
`define T_clk 10
module mux()
// main testbench related parameters 
`define INSTRUCTIONS_FILE "/home/matteo/git/RV-MAGIC/main/tb/hex_mc/fwd_load_alu.riscv"
`define RANDOM_DATA_FILE "../../main/tb/hex_mc/dmemh.mem"
`define NUMBER_OF_INSTRUCTIONS 10

// clock period
`define T_clk 10
// main testbench related parameters 
`define INSTRUCTIONS_FILE "../../main/tb/mc/1-instr_list_no_jump.riscv"
`define RANDOM_DATA_FILE "../../main/tb/mc/3-fwd_test.riscv"
`define NUMBER_OF_INSTRUCTIONS 10

// clock period
`define T_clk 20
`define half_T_clk 10
// main testbench related parameters 
`define INSTRUCTIONS_FILE "../../main/tb/hex_mc/2-instr_list_w_jumps.mc.riscv"
`define RANDOM_DATA_FILE "../../main/tb/hex_mc/3-fwd_test.mc.riscv"
`define NUMBER_OF_INSTRUCTIONS 10

// clock period
`define T_clk 4
// main testbench related parameters 
`define INSTRUCTIONS_FILE "../../main/tb/instructions.txt"
`define RANDOM_DATA_FILE "../../main/tb/random_data.txt"
`define NUMBER_OF_INSTRUCTIONS 10

`define T_clk 20
// width-related constants
`define INST_WIDTH      32
`define ADDR_WIDTH      32
`define WORD_WIDTH      32
`define HWORD_WIDTH     16
`define BYTE_WIDTH      8
`define SHAMT_WIDTH     5
`define RF_ADDR_WIDTH   5

// U-type opcodes
`define RV32_LUI     7'b0110111
`define RV32_AUIPC   7'b0010111

// J-type opcodes
`define RV32_JAL     7'b1101111

// I-type opcodes
`define RV32_JALR    7'b1100111
`define RV32_LOAD    7'b0000011
`define RV32_OP_IMM  7'b0010011
`define RV32_FENCE   7'b0001111
`define RV32_SYSTEM  7'b1110011

// B-type opcodes
`define RV32_BRANCH  7'b1100011

// S-type opcodes
`define RV32_STORE   7'b0100011

// R-type opcodes
`define RV32_OP      7'b0110011

// NOP
`define RV_NOP `INST_WIDTH'b0010011

// arithmetic funct3 encodings
`define FUNCT3_ADD_SUB 0
`define FUNCT3_SLL     1
`define FUNCT3_SLT     2
`define FUNCT3_SLTU    3
`define FUNCT3_XOR     4
`define FUNCT3_SRA_SRL 5
`define FUNCT3_OR      6
`define FUNCT3_AND     7

// branch funct3 encodings
`define FUNCT3_BEQ  0
`define FUNCT3_BNE  1
`define FUNCT3_BLT  4
`define FUNCT3_BGE  5
`define FUNCT3_BLTU 6
`define FUNCT3_BGEU 7

// fence funct3 encodings
`define FUNCT3_FENCE   0
`define FUNCT3_FENCE_I 1

// system funct3 encodings
`define FUNCT3_ENV    0
`define FUNCT3_CSRRW  1
`define FUNCT3_CSRRS  2
`define FUNCT3_CSRRC  3
`define FUNCT3_CSRRWI 5
`define FUNCT3_CSRRSI 6
`define FUNCT3_CSRRCI 7

// env funct12 encodings
`define FUNCT12_ECALL  12'b000000000000
`define FUNCT12_EBREAK 12'b000000000001













// width for MUX control inside immediate generation

`define IMMEDIATE_SELECTION_WIDTH 3

// widths
`define RV32I_OPCODE_WIDTH  7
`define RV32I_FUNCT3_WIDTH 3
`define RV32I_SHAMT_WIDTH 5
`define RV32I_FUNCT7_WIDTH 7

// instruction types

`define R_TYPE `IMMEDIATE_SELECTION_WIDTH'b101
`define I_TYPE `IMMEDIATE_SELECTION_WIDTH'b000
`define S_TYPE `IMMEDIATE_SELECTION_WIDTH'b001
`define B_TYPE `IMMEDIATE_SELECTION_WIDTH'b010
`define U_TYPE `IMMEDIATE_SELECTION_WIDTH'b011
`define J_TYPE `IMMEDIATE_SELECTION_WIDTH'b100

// bit positions
`define RV32I_FUNCT7_START 25
`define RV32I_OPCODE_START 0
`define RV32I_FUNCT3_START 12
`define RV32I_SHAMT_START 20


// operations
`define RV32I_LUI_OPCODE `RV32I_OPCODE_WIDTH'b0110111 // U-type
`define RV32I_AUIPC_OPCODE `RV32I_OPCODE_WIDTH'b0010111 // U-type
`define RV32I_JAL_OPCODE `RV32I_OPCODE_WIDTH'b1101111 // J-type
`define RV32I_JALR_OPCODE `RV32I_OPCODE_WIDTH'b1100111 // I-type
`define RV32I_BEQ_OPCODE `RV32I_OPCODE_WIDTH'b1100011 // B-type
`define RV32I_BNE_OPCODE `RV32I_OPCODE_WIDTH'b1100011 // B-type
`define RV32I_BLT_OPCODE `RV32I_OPCODE_WIDTH'b1100011 // B-type
`define RV32I_BGE_OPCODE `RV32I_OPCODE_WIDTH'b1100011 // B-type
`define RV32I_BLTU_OPCODE `RV32I_OPCODE_WIDTH'b1100011 // B-type
`define RV32I_BGEU_OPCODE `RV32I_OPCODE_WIDTH'b1100011 // B-type
`define RV32I_LB_OPCODE `RV32I_OPCODE_WIDTH'b0000011 // I-type
`define RV32I_LH_OPCODE `RV32I_OPCODE_WIDTH'b0000011 // I-type
`define RV32I_LW_OPCODE `RV32I_OPCODE_WIDTH'b0000011 // I-type
`define RV32I_LBU_OPCODE `RV32I_OPCODE_WIDTH'b0000011 // I-type
`define RV32I_LHU_OPCODE `RV32I_OPCODE_WIDTH'b0000011 // I-type
`define RV32I_SB_OPCODE `RV32I_OPCODE_WIDTH'b0100011 // S-type
`define RV32I_SH_OPCODE `RV32I_OPCODE_WIDTH'b0100011 // S-type
`define RV32I_SW_OPCODE `RV32I_OPCODE_WIDTH'b0100011 // S-type
`define RV32I_ADDI_OPCODE `RV32I_OPCODE_WIDTH'b0010011 // I-type
`define RV32I_SLTI_OPCODE `RV32I_OPCODE_WIDTH'b0010011 // I-type
`define RV32I_SLTIU_OPCODE `RV32I_OPCODE_WIDTH'b0010011 // I-type
`define RV32I_XORI_OPCODE `RV32I_OPCODE_WIDTH'b0010011 // I-type
`define RV32I_ORI_OPCODE `RV32I_OPCODE_WIDTH'b0010011 // I-type
`define RV32I_ANDI_OPCODE `RV32I_OPCODE_WIDTH'b0010011 // I-type
`define RV32I_SLLI_OPCODE `RV32I_OPCODE_WIDTH'b0010011 // R-type
`define RV32I_SRLI_OPCODE `RV32I_OPCODE_WIDTH'b0010011 // R-type
`define RV32I_SRAI_OPCODE `RV32I_OPCODE_WIDTH'b0010011 // R-type
`define RV32I_ADD_OPCODE `RV32I_OPCODE_WIDTH'b0110011 // R-type
`define RV32I_SUB_OPCODE `RV32I_OPCODE_WIDTH'b0110011 // R-type
`define RV32I_SLL_OPCODE `RV32I_OPCODE_WIDTH'b0110011 // R-type
`define RV32I_SLT_OPCODE `RV32I_OPCODE_WIDTH'b0110011 // R-type
`define RV32I_SLTU_OPCODE `RV32I_OPCODE_WIDTH'b0110011 // R-type
`define RV32I_XOR_OPCODE `RV32I_OPCODE_WIDTH'b0110011 // R-type
`define RV32I_SRL_OPCODE `RV32I_OPCODE_WIDTH'b0110011 // R-type
`define RV32I_SRA_OPCODE `RV32I_OPCODE_WIDTH'b0110011 // R-type
`define RV32I_OR_OPCODE `RV32I_OPCODE_WIDTH'b0110011 // R-type
`define RV32I_AND_OPCODE `RV32I_OPCODE_WIDTH'b0110011 // R-type
// FOLLOWING INSTRUCTIONS ARE DEFINED BUT NOT USED
`define RV32I_FENCE_OPCODE `RV32I_OPCODE_WIDTH'b0001111
`define RV32I_FENCE_I_OPCODE `RV32I_OPCODE_WIDTH'b0001111
`define RV32I_ECALL_OPCODE `RV32I_OPCODE_WIDTH'b1110011
`define RV32I_EBREAK_OPCODE `RV32I_OPCODE_WIDTH'b1110011
`define RV32I_CSRRW_OPCODE `RV32I_OPCODE_WIDTH'b1110011
`define RV32I_CSRRS_OPCODE `RV32I_OPCODE_WIDTH'b1110011
`define RV32I_CSRRC_OPCODE `RV32I_OPCODE_WIDTH'b1110011
`define RV32I_CSRRWI_OPCODE `RV32I_OPCODE_WIDTH'b1110011
`define RV32I_CSRRSI_OPCODE `RV32I_OPCODE_WIDTH'b1110011
`define RV32I_CSRRCI_OPCODE `RV32I_OPCODE_WIDTH'b1110011


// funct3 codes
`define RV32I_JALR_FUNCT3 `RV32I_FUNCT3_WIDTH'b000
`define RV32I_BEQ_FUNCT3 `RV32I_FUNCT3_WIDTH'b000
`define RV32I_BNE_FUNCT3 `RV32I_FUNCT3_WIDTH'b001
`define RV32I_BLT_FUNCT3 `RV32I_FUNCT3_WIDTH'b100
`define RV32I_BGE_FUNCT3 `RV32I_FUNCT3_WIDTH'b101
`define RV32I_BLTU_FUNCT3 `RV32I_FUNCT3_WIDTH'b110
`define RV32I_BGEU_FUNCT3 `RV32I_FUNCT3_WIDTH'b111
`define RV32I_LB_FUNCT3 `RV32I_FUNCT3_WIDTH'b000
`define RV32I_LH_FUNCT3 `RV32I_FUNCT3_WIDTH'b001
`define RV32I_LW_FUNCT3 `RV32I_FUNCT3_WIDTH'b010
`define RV32I_LBU_FUNCT3 `RV32I_FUNCT3_WIDTH'b100
`define RV32I_LHU_FUNCT3 `RV32I_FUNCT3_WIDTH'b101
`define RV32I_SB_FUNCT3 `RV32I_FUNCT3_WIDTH'b000
`define RV32I_SH_FUNCT3 `RV32I_FUNCT3_WIDTH'b001
`define RV32I_SW_FUNCT3 `RV32I_FUNCT3_WIDTH'b010
`define RV32I_ADDI_FUNCT3 `RV32I_FUNCT3_WIDTH'b000
`define RV32I_SLTI_FUNCT3 `RV32I_FUNCT3_WIDTH'b010
`define RV32I_SLTIU_FUNCT3 `RV32I_FUNCT3_WIDTH'b011
`define RV32I_XORI_FUNCT3 `RV32I_FUNCT3_WIDTH'b100
`define RV32I_ORI_FUNCT3 `RV32I_FUNCT3_WIDTH'b110
`define RV32I_ANDI_FUNCT3 `RV32I_FUNCT3_WIDTH'b111
`define RV32I_SLLI_FUNCT3 `RV32I_FUNCT3_WIDTH'b001
`define RV32I_SRLI_FUNCT3 `RV32I_FUNCT3_WIDTH'b101
`define RV32I_SRAI_FUNCT3 `RV32I_FUNCT3_WIDTH'b101
`define RV32I_ADD_FUNCT3 `RV32I_FUNCT3_WIDTH'b000
`define RV32I_SUB_FUNCT3 `RV32I_FUNCT3_WIDTH'b000
`define RV32I_SLL_FUNCT3 `RV32I_FUNCT3_WIDTH'b001
`define RV32I_SLT_FUNCT3 `RV32I_FUNCT3_WIDTH'b010
`define RV32I_SLTU_FUNCT3 `RV32I_FUNCT3_WIDTH'b011
`define RV32I_XOR_FUNCT3 `RV32I_FUNCT3_WIDTH'b100
`define RV32I_SRL_FUNCT3 `RV32I_FUNCT3_WIDTH'b101
`define RV32I_SRA_FUNCT3 `RV32I_FUNCT3_WIDTH'b101
`define RV32I_OR_FUNCT3 `RV32I_FUNCT3_WIDTH'b110
`define RV32I_AND_FUNCT3 `RV32I_FUNCT3_WIDTH'b111
// FOLLOWING INSTRUCTIONS ARE DEFINED BUT NOT USED
`define RV32I_FENCE_FUNCT3 `RV32I_FUNCT3_WIDTH'b000
`define RV32I_FENCE_I_FUNCT3 `RV32I_FUNCT3_WIDTH'b001
`define RV32I_ECALL_FUNCT3 `RV32I_FUNCT3_WIDTH'b000
`define RV32I_EBREAK_FUNCT3 `RV32I_FUNCT3_WIDTH'b000
`define RV32I_CSRRW_FUNCT3 `RV32I_FUNCT3_WIDTH'b001
`define RV32I_CSRRS_FUNCT3 `RV32I_FUNCT3_WIDTH'b010
`define RV32I_CSRRC_FUNCT3 `RV32I_FUNCT3_WIDTH'b011
`define RV32I_CSRRWI_FUNCT3 `RV32I_FUNCT3_WIDTH'b101
`define RV32I_CSRRSI_FUNCT3 `RV32I_FUNCT3_WIDTH'b110
`define RV32I_CSRRCI_FUNCT3 `RV32I_FUNCT3_WIDTH'b111


// funct7 codes
`define RV32I_SLLI_FUNCT7 `RV32I_FUNCT7_WIDTH'b0000000
`define RV32I_SRLI_FUNCT7 `RV32I_FUNCT7_WIDTH'b0000000
`define RV32I_SRAI_FUNCT7 `RV32I_FUNCT7_WIDTH'b0100000
`define RV32I_ADD_FUNCT7 `RV32I_FUNCT7_WIDTH'b0000000
`define RV32I_SUB_FUNCT7 `RV32I_FUNCT7_WIDTH'b0100000
`define RV32I_SLL_FUNCT7 `RV32I_FUNCT7_WIDTH'b0000000
`define RV32I_SLT_FUNCT7 `RV32I_FUNCT7_WIDTH'b0000000
`define RV32I_SLTU_FUNCT7 `RV32I_FUNCT7_WIDTH'b0000000
`define RV32I_XOR_FUNCT7 `RV32I_FUNCT7_WIDTH'b0000000
`define RV32I_SRL_FUNCT7 `RV32I_FUNCT7_WIDTH'b0000000
`define RV32I_SRA_FUNCT7 `RV32I_FUNCT7_WIDTH'b0100000
`define RV32I_OR_FUNCT7 `RV32I_FUNCT7_WIDTH'b0000000
`define RV32I_AND_FUNCT7 `RV32I_FUNCT7_WIDTH'b0000000

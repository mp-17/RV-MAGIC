// main testbench related parameters 
`define INSTRUCTIONS_FILE "/home/michi/Documents/git-projects/RV-MAGIC/main/tb/hex_mc/ass_test.riscv"
`define RANDOM_DATA_FILE "../../main/tb/hex_mc/dmemh.mem"
`define NUMBER_OF_INSTRUCTIONS 10

// clock period
`define T_clk 10